`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/11/25 16:47:49
// Design Name: 
// Module Name: ALU
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module Adder(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
    );
    assign sum[0] = a[0] ^ b[0] ^ 0;
    assign sum[1] = a[1] ^ b[1] ^ (a[0] * b[0] + (a[0] ^ b[0]) * 0);
    assign sum[2] = a[2] ^ b[2] ^ (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0));
    assign sum[3] = a[3] ^ b[3] ^ (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)));
    assign sum[4] = a[4] ^ b[4] ^ (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))));
    assign sum[5] = a[5] ^ b[5] ^ (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))));
    assign sum[6] = a[6] ^ b[6] ^ (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))));
    assign sum[7] = a[7] ^ b[7] ^ (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))));
    assign sum[8] = a[8] ^ b[8] ^ (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))));
    assign sum[9] = a[9] ^ b[9] ^ (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))));
    assign sum[10] = a[10] ^ b[10] ^ (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))));
    assign sum[11] = a[11] ^ b[11] ^ (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))));
    assign sum[12] = a[12] ^ b[12] ^ (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))));
    assign sum[13] = a[13] ^ b[13] ^ (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))));
    assign sum[14] = a[14] ^ b[14] ^ (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))));
    assign sum[15] = a[15] ^ b[15] ^ (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))));
    assign sum[16] = a[16] ^ b[16] ^ (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))));
    assign sum[17] = a[17] ^ b[17] ^ (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))));
    assign sum[18] = a[18] ^ b[18] ^ (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))));
    assign sum[19] = a[19] ^ b[19] ^ (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))));
    assign sum[20] = a[20] ^ b[20] ^ (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))));
    assign sum[21] = a[21] ^ b[21] ^ (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))));
    assign sum[22] = a[22] ^ b[22] ^ (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))));
    assign sum[23] = a[23] ^ b[23] ^ (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))));
    assign sum[24] = a[24] ^ b[24] ^ (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))))));
    assign sum[25] = a[25] ^ b[25] ^ (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))))));
    assign sum[26] = a[26] ^ b[26] ^ (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))))))));
    assign sum[27] = a[27] ^ b[27] ^ (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))))))));
    assign sum[28] = a[28] ^ b[28] ^ (a[27] * b[27] + (a[27] ^ b[27]) * (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))))))))));
    assign sum[29] = a[29] ^ b[29] ^ (a[28] * b[28] + (a[28] ^ b[28]) * (a[27] * b[27] + (a[27] ^ b[27]) * (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))))))))));
    assign sum[30] = a[30] ^ b[30] ^ (a[29] * b[29] + (a[29] ^ b[29]) * (a[28] * b[28] + (a[28] ^ b[28]) * (a[27] * b[27] + (a[27] ^ b[27]) * (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))))))))))));
    assign sum[31] = a[31] ^ b[31] ^ (a[30] * b[30] + (a[30] ^ b[30]) * (a[29] * b[29] + (a[29] ^ b[29]) * (a[28] * b[28] + (a[28] ^ b[28]) * (a[27] * b[27] + (a[27] ^ b[27]) * (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))))))))))));
endmodule

module Shift(input [31:0] B, input[3:0] Op, input [31:0] A, input usigned,output [31:0] res);
	wire [31:0] left_shift;
	wire [31:0] right_shift;
	wire [31:0] aright_shift;

	assign left_shift = B << A;
	assign right_shift = B >> A;
	assign aright_shift = $signed(B)>>> A;

	assign res = (Op[0] == 1)? left_shift : (usigned == 1? aright_shift : right_shift);
endmodule

module BitOp(input[31:0] A, input[31:0] B, input[3:0] Op, output [31:0] res);
	wire [31:0] and_res;
	wire [31:0] or_res;
	wire [31:0] xor_res;
	wire [31:0] nor_res;
	
	assign and_res = A & B;
	assign or_res = A | B;
	assign xor_res = A ^ B;
	assign nor_res = ~or_res;

	assign res = Op[2] == 0? (Op[0] == 0? and_res : or_res) : (Op[0] == 0 ? xor_res : nor_res);
endmodule

module Leg(input[31:0] A, input[31:0] B, input[3:0] Op ,input usigned,output [31:0] res);
    wire less_res, less_equal_res;
    wire greater_res, greater_equal_res;
    wire less_v_res, unsigned_less_v_res, unsigned_less_res;
    wire eq_res;
    
	assign less_v_res = $signed(A) < $signed(B);
	assign unsigned_less_v_res = A < B;
    assign less_res = $signed(A) < 0;  
	assign less_equal_res = $signed(A) <= 0;
	assign greater_equal_res = $signed(A) >= 0;
	assign greater_res = $signed(A) > 0;
	assign eq_res = A == B;
	
	assign res = (~Op[3]&&~Op[2]&&~Op[1])?eq_res:(Op[2]==0 && Op[1]==0 && Op[0]==1) ? (usigned==1 ? unsigned_less_v_res: less_v_res):(Op[2]==1 ? (Op[0]==1 ? greater_equal_res : less_res):(Op[0]==1 ? greater_res : less_equal_res)); 	
endmodule

 module ALU(PC, PCSrc, A, B, Op, usigned, C, zero, over);
    input [31:0] PC;
    input [31:0] A;
    input [31:0] B;
    input [3:0] Op;
    input [2:0] PCSrc;
    input usigned;
    output [31:0] C;
    output zero;
    output over;
    
    wire [31:0] shift_res, aoxn_res, sum_res, leg_res, PC_res;
    wire [31:0] neg_B, b_input;
	wire cout;
	Adder neg(~B, 32'b1, neg_B);
	assign b_input = Op[0]? neg_B : B;
    
    Shift shift(B, Op, A, usigned, shift_res);
	BitOp bitOp(A, B, Op, aoxn_res);
	Adder adder(A, b_input, sum_res);
	Adder adder_pc(PC, 32'b1000, PC_res);
    Leg leg(A, B, Op, usigned, leg_res);
    
	assign over = (~Op[3] & ~Op[2] & ~Op[1]) ? ((usigned) & ((A[31] == b_input[31]) & (A[31] != sum_res[31]))) : 0;
    
    assign C = (PCSrc == 3'b011)? PC_res : (Op[3]? ((~Op[2] & ~Op[1] & Op[0])? leg_res : shift_res) : ((~Op[2] & ~Op[1])? sum_res : (Op[2] & Op[1])? (B << 16) : aoxn_res));
    
    assign zero = (C == 0) ? 1 : 0;
endmodule

