`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/11/03 16:23:57
// Design Name: 
// Module Name: Adder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Adder(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
    );
    assign sum[0] = a[0] ^ b[0] ^ 0;
    assign sum[1] = a[1] ^ b[1] ^ (a[0] * b[0] + (a[0] ^ b[0]) * 0);
    assign sum[2] = a[2] ^ b[2] ^ (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0));
    assign sum[3] = a[3] ^ b[3] ^ (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)));
    assign sum[4] = a[4] ^ b[4] ^ (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))));
    assign sum[5] = a[5] ^ b[5] ^ (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))));
    assign sum[6] = a[6] ^ b[6] ^ (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))));
    assign sum[7] = a[7] ^ b[7] ^ (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))));
    assign sum[8] = a[8] ^ b[8] ^ (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))));
    assign sum[9] = a[9] ^ b[9] ^ (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))));
    assign sum[10] = a[10] ^ b[10] ^ (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))));
    assign sum[11] = a[11] ^ b[11] ^ (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))));
    assign sum[12] = a[12] ^ b[12] ^ (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))));
    assign sum[13] = a[13] ^ b[13] ^ (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))));
    assign sum[14] = a[14] ^ b[14] ^ (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))));
    assign sum[15] = a[15] ^ b[15] ^ (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))));
    assign sum[16] = a[16] ^ b[16] ^ (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))));
    assign sum[17] = a[17] ^ b[17] ^ (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))));
    assign sum[18] = a[18] ^ b[18] ^ (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))));
    assign sum[19] = a[19] ^ b[19] ^ (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))));
    assign sum[20] = a[20] ^ b[20] ^ (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))));
    assign sum[21] = a[21] ^ b[21] ^ (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))));
    assign sum[22] = a[22] ^ b[22] ^ (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))));
    assign sum[23] = a[23] ^ b[23] ^ (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))));
    assign sum[24] = a[24] ^ b[24] ^ (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))))));
    assign sum[25] = a[25] ^ b[25] ^ (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))))));
    assign sum[26] = a[26] ^ b[26] ^ (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))))))));
    assign sum[27] = a[27] ^ b[27] ^ (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))))))));
    assign sum[28] = a[28] ^ b[28] ^ (a[27] * b[27] + (a[27] ^ b[27]) * (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))))))))));
    assign sum[29] = a[29] ^ b[29] ^ (a[28] * b[28] + (a[28] ^ b[28]) * (a[27] * b[27] + (a[27] ^ b[27]) * (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))))))))));
    assign sum[30] = a[30] ^ b[30] ^ (a[29] * b[29] + (a[29] ^ b[29]) * (a[28] * b[28] + (a[28] ^ b[28]) * (a[27] * b[27] + (a[27] ^ b[27]) * (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0))))))))))))))))))))))))))))));
    assign sum[31] = a[31] ^ b[31] ^ (a[30] * b[30] + (a[30] ^ b[30]) * (a[29] * b[29] + (a[29] ^ b[29]) * (a[28] * b[28] + (a[28] ^ b[28]) * (a[27] * b[27] + (a[27] ^ b[27]) * (a[26] * b[26] + (a[26] ^ b[26]) * (a[25] * b[25] + (a[25] ^ b[25]) * (a[24] * b[24] + (a[24] ^ b[24]) * (a[23] * b[23] + (a[23] ^ b[23]) * (a[22] * b[22] + (a[22] ^ b[22]) * (a[21] * b[21] + (a[21] ^ b[21]) * (a[20] * b[20] + (a[20] ^ b[20]) * (a[19] * b[19] + (a[19] ^ b[19]) * (a[18] * b[18] + (a[18] ^ b[18]) * (a[17] * b[17] + (a[17] ^ b[17]) * (a[16] * b[16] + (a[16] ^ b[16]) * (a[15] * b[15] + (a[15] ^ b[15]) * (a[14] * b[14] + (a[14] ^ b[14]) * (a[13] * b[13] + (a[13] ^ b[13]) * (a[12] * b[12] + (a[12] ^ b[12]) * (a[11] * b[11] + (a[11] ^ b[11]) * (a[10] * b[10] + (a[10] ^ b[10]) * (a[9] * b[9] + (a[9] ^ b[9]) * (a[8] * b[8] + (a[8] ^ b[8]) * (a[7] * b[7] + (a[7] ^ b[7]) * (a[6] * b[6] + (a[6] ^ b[6]) * (a[5] * b[5] + (a[5] ^ b[5]) * (a[4] * b[4] + (a[4] ^ b[4]) * (a[3] * b[3] + (a[3] ^ b[3]) * (a[2] * b[2] + (a[2] ^ b[2]) * (a[1] * b[1] + (a[1] ^ b[1]) * (a[0] * b[0] + (a[0] ^ b[0]) * 0)))))))))))))))))))))))))))))));
endmodule
